// i2c_controller.sv - Reed Foster
// controller for ADAU1761 control interface

module i2c_controller (
  input wire clk, reset,
  output  scl,
  input   sda_i,
  output  sda_o,
  output  sda_t
);

enum {


endmodule
